`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2017/11/02 14:44:10
// Design Name: 
// Module Name: mux2
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module mux2 #(
	parameter 					WIDTH = 8
)(
	input		[WIDTH-1:0] 	din0,
	input		[WIDTH-1:0] 	din1,
	input						sel_i,
	output 		[WIDTH-1:0] 	dout
    );
	//add your code here
	assign dout = sel_i ? din1 : din0;
endmodule
